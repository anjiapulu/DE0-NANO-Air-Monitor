// DE0_NANO_QSYS.v

// Generated using ACDS version 13.1 162 at 2021.07.30.14:26:14

`timescale 1 ps / 1 ps
module DE0_NANO_QSYS (
		input  wire        clk_clk,                             //                             clk.clk
		input  wire        reset_reset_n,                       //                           reset.reset_n
		input  wire        key_external_connection_export,      //         key_external_connection.export
		output wire [12:0] sdram_wire_addr,                     //                      sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                       //                                .ba
		output wire        sdram_wire_cas_n,                    //                                .cas_n
		output wire        sdram_wire_cke,                      //                                .cke
		output wire        sdram_wire_cs_n,                     //                                .cs_n
		inout  wire [15:0] sdram_wire_dq,                       //                                .dq
		output wire [1:0]  sdram_wire_dqm,                      //                                .dqm
		output wire        sdram_wire_ras_n,                    //                                .ras_n
		output wire        sdram_wire_we_n,                     //                                .we_n
		output wire        altpll_sdram_clk,                    //                    altpll_sdram.clk
		input  wire        altpll_areset_conduit_export,        //           altpll_areset_conduit.export
		output wire        altpll_locked_conduit_export,        //           altpll_locked_conduit.export
		output wire        altpll_phasedone_conduit_export,     //        altpll_phasedone_conduit.export
		output wire        scl_export,                          //                             scl.export
		inout  wire        sda_export,                          //                             sda.export
		input  wire        uart_test_external_connection_rxd,   //   uart_test_external_connection.rxd
		output wire        uart_test_external_connection_txd,   //                                .txd
		input  wire        uart_co_external_connection_rxd,     //     uart_co_external_connection.rxd
		output wire        uart_co_external_connection_txd,     //                                .txd
		input  wire        uart_sds011_external_connection_rxd, // uart_sds011_external_connection.rxd
		output wire        uart_sds011_external_connection_txd, //                                .txd
		input  wire        uart_so2_external_connection_rxd,    //    uart_so2_external_connection.rxd
		output wire        uart_so2_external_connection_txd,    //                                .txd
		input  wire        uart_o3_external_connection_rxd,     //     uart_o3_external_connection.rxd
		output wire        uart_o3_external_connection_txd,     //                                .txd
		input  wire        uart_hmi_external_connection_rxd,    //    uart_hmi_external_connection.rxd
		output wire        uart_hmi_external_connection_txd,    //                                .txd
		output wire        epcs_flash_external_dclk,            //             epcs_flash_external.dclk
		output wire        epcs_flash_external_sce,             //                                .sce
		output wire        epcs_flash_external_sdo,             //                                .sdo
		input  wire        epcs_flash_external_data0            //                                .data0
	);

	wire         altpll_c0_clk;                                              // altpll:c0 -> [irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, irq_synchronizer_002:sender_clk, irq_synchronizer_003:sender_clk, irq_synchronizer_004:sender_clk, irq_synchronizer_005:sender_clk, irq_synchronizer_006:sender_clk, jtag_uart:clk, key:clk, mm_interconnect_0:altpll_c0_clk, nios2_qsys:clk, rst_controller:clk, sdram:clk, sysid_qsys:clock]
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                         // mm_interconnect_0:key_s1_writedata -> key:writedata
	wire   [1:0] mm_interconnect_0_key_s1_address;                           // mm_interconnect_0:key_s1_address -> key:address
	wire         mm_interconnect_0_key_s1_chipselect;                        // mm_interconnect_0:key_s1_chipselect -> key:chipselect
	wire         mm_interconnect_0_key_s1_write;                             // mm_interconnect_0:key_s1_write -> key:write_n
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                          // key:readdata -> mm_interconnect_0:key_s1_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest; // nios2_qsys:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_jtag_debug_module_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_jtag_debug_module_address -> nios2_qsys:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_jtag_debug_module_write -> nios2_qsys:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_jtag_debug_module_read -> nios2_qsys:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata;    // nios2_qsys:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_jtag_debug_module_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_jtag_debug_module_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_writedata;   // mm_interconnect_0:epcs_flash_epcs_control_port_writedata -> epcs_flash:writedata
	wire   [8:0] mm_interconnect_0_epcs_flash_epcs_control_port_address;     // mm_interconnect_0:epcs_flash_epcs_control_port_address -> epcs_flash:address
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_chipselect;  // mm_interconnect_0:epcs_flash_epcs_control_port_chipselect -> epcs_flash:chipselect
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_write;       // mm_interconnect_0:epcs_flash_epcs_control_port_write -> epcs_flash:write_n
	wire         mm_interconnect_0_epcs_flash_epcs_control_port_read;        // mm_interconnect_0:epcs_flash_epcs_control_port_read -> epcs_flash:read_n
	wire  [31:0] mm_interconnect_0_epcs_flash_epcs_control_port_readdata;    // epcs_flash:readdata -> mm_interconnect_0:epcs_flash_epcs_control_port_readdata
	wire  [15:0] mm_interconnect_0_uart_sds011_s1_writedata;                 // mm_interconnect_0:uart_sds011_s1_writedata -> uart_sds011:writedata
	wire   [2:0] mm_interconnect_0_uart_sds011_s1_address;                   // mm_interconnect_0:uart_sds011_s1_address -> uart_sds011:address
	wire         mm_interconnect_0_uart_sds011_s1_chipselect;                // mm_interconnect_0:uart_sds011_s1_chipselect -> uart_sds011:chipselect
	wire         mm_interconnect_0_uart_sds011_s1_write;                     // mm_interconnect_0:uart_sds011_s1_write -> uart_sds011:write_n
	wire         mm_interconnect_0_uart_sds011_s1_read;                      // mm_interconnect_0:uart_sds011_s1_read -> uart_sds011:read_n
	wire  [15:0] mm_interconnect_0_uart_sds011_s1_readdata;                  // uart_sds011:readdata -> mm_interconnect_0:uart_sds011_s1_readdata
	wire         mm_interconnect_0_uart_sds011_s1_begintransfer;             // mm_interconnect_0:uart_sds011_s1_begintransfer -> uart_sds011:begintransfer
	wire         nios2_qsys_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_data_master_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                           // nios2_qsys:d_writedata -> mm_interconnect_0:nios2_qsys_data_master_writedata
	wire  [25:0] nios2_qsys_data_master_address;                             // nios2_qsys:d_address -> mm_interconnect_0:nios2_qsys_data_master_address
	wire         nios2_qsys_data_master_write;                               // nios2_qsys:d_write -> mm_interconnect_0:nios2_qsys_data_master_write
	wire         nios2_qsys_data_master_read;                                // nios2_qsys:d_read -> mm_interconnect_0:nios2_qsys_data_master_read
	wire  [31:0] nios2_qsys_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_data_master_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                         // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_data_master_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_data_master_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                          // nios2_qsys:d_byteenable -> mm_interconnect_0:nios2_qsys_data_master_byteenable
	wire  [31:0] mm_interconnect_0_scl_s1_writedata;                         // mm_interconnect_0:scl_s1_writedata -> scl:writedata
	wire   [1:0] mm_interconnect_0_scl_s1_address;                           // mm_interconnect_0:scl_s1_address -> scl:address
	wire         mm_interconnect_0_scl_s1_chipselect;                        // mm_interconnect_0:scl_s1_chipselect -> scl:chipselect
	wire         mm_interconnect_0_scl_s1_write;                             // mm_interconnect_0:scl_s1_write -> scl:write_n
	wire  [31:0] mm_interconnect_0_scl_s1_readdata;                          // scl:readdata -> mm_interconnect_0:scl_s1_readdata
	wire  [31:0] mm_interconnect_0_sda_s1_writedata;                         // mm_interconnect_0:sda_s1_writedata -> sda:writedata
	wire   [1:0] mm_interconnect_0_sda_s1_address;                           // mm_interconnect_0:sda_s1_address -> sda:address
	wire         mm_interconnect_0_sda_s1_chipselect;                        // mm_interconnect_0:sda_s1_chipselect -> sda:chipselect
	wire         mm_interconnect_0_sda_s1_write;                             // mm_interconnect_0:sda_s1_write -> sda:write_n
	wire  [31:0] mm_interconnect_0_sda_s1_readdata;                          // sda:readdata -> mm_interconnect_0:sda_s1_readdata
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_writedata;               // mm_interconnect_0:altpll_pll_slave_writedata -> altpll:writedata
	wire   [1:0] mm_interconnect_0_altpll_pll_slave_address;                 // mm_interconnect_0:altpll_pll_slave_address -> altpll:address
	wire         mm_interconnect_0_altpll_pll_slave_write;                   // mm_interconnect_0:altpll_pll_slave_write -> altpll:write
	wire         mm_interconnect_0_altpll_pll_slave_read;                    // mm_interconnect_0:altpll_pll_slave_read -> altpll:read
	wire  [31:0] mm_interconnect_0_altpll_pll_slave_readdata;                // altpll:readdata -> mm_interconnect_0:altpll_pll_slave_readdata
	wire  [15:0] mm_interconnect_0_uart_no2_s1_writedata;                    // mm_interconnect_0:uart_no2_s1_writedata -> uart_no2:writedata
	wire   [2:0] mm_interconnect_0_uart_no2_s1_address;                      // mm_interconnect_0:uart_no2_s1_address -> uart_no2:address
	wire         mm_interconnect_0_uart_no2_s1_chipselect;                   // mm_interconnect_0:uart_no2_s1_chipselect -> uart_no2:chipselect
	wire         mm_interconnect_0_uart_no2_s1_write;                        // mm_interconnect_0:uart_no2_s1_write -> uart_no2:write_n
	wire         mm_interconnect_0_uart_no2_s1_read;                         // mm_interconnect_0:uart_no2_s1_read -> uart_no2:read_n
	wire  [15:0] mm_interconnect_0_uart_no2_s1_readdata;                     // uart_no2:readdata -> mm_interconnect_0:uart_no2_s1_readdata
	wire         mm_interconnect_0_uart_no2_s1_begintransfer;                // mm_interconnect_0:uart_no2_s1_begintransfer -> uart_no2:begintransfer
	wire         nios2_qsys_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_instruction_master_waitrequest -> nios2_qsys:i_waitrequest
	wire  [25:0] nios2_qsys_instruction_master_address;                      // nios2_qsys:i_address -> mm_interconnect_0:nios2_qsys_instruction_master_address
	wire         nios2_qsys_instruction_master_read;                         // nios2_qsys:i_read -> mm_interconnect_0:nios2_qsys_instruction_master_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_instruction_master_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_instruction_master_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                     // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                       // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                         // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                      // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                           // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                            // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                        // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                   // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                      // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [15:0] mm_interconnect_0_uart_co_s1_writedata;                     // mm_interconnect_0:uart_co_s1_writedata -> uart_co:writedata
	wire   [2:0] mm_interconnect_0_uart_co_s1_address;                       // mm_interconnect_0:uart_co_s1_address -> uart_co:address
	wire         mm_interconnect_0_uart_co_s1_chipselect;                    // mm_interconnect_0:uart_co_s1_chipselect -> uart_co:chipselect
	wire         mm_interconnect_0_uart_co_s1_write;                         // mm_interconnect_0:uart_co_s1_write -> uart_co:write_n
	wire         mm_interconnect_0_uart_co_s1_read;                          // mm_interconnect_0:uart_co_s1_read -> uart_co:read_n
	wire  [15:0] mm_interconnect_0_uart_co_s1_readdata;                      // uart_co:readdata -> mm_interconnect_0:uart_co_s1_readdata
	wire         mm_interconnect_0_uart_co_s1_begintransfer;                 // mm_interconnect_0:uart_co_s1_begintransfer -> uart_co:begintransfer
	wire  [15:0] mm_interconnect_0_uart_so2_s1_writedata;                    // mm_interconnect_0:uart_so2_s1_writedata -> uart_so2:writedata
	wire   [2:0] mm_interconnect_0_uart_so2_s1_address;                      // mm_interconnect_0:uart_so2_s1_address -> uart_so2:address
	wire         mm_interconnect_0_uart_so2_s1_chipselect;                   // mm_interconnect_0:uart_so2_s1_chipselect -> uart_so2:chipselect
	wire         mm_interconnect_0_uart_so2_s1_write;                        // mm_interconnect_0:uart_so2_s1_write -> uart_so2:write_n
	wire         mm_interconnect_0_uart_so2_s1_read;                         // mm_interconnect_0:uart_so2_s1_read -> uart_so2:read_n
	wire  [15:0] mm_interconnect_0_uart_so2_s1_readdata;                     // uart_so2:readdata -> mm_interconnect_0:uart_so2_s1_readdata
	wire         mm_interconnect_0_uart_so2_s1_begintransfer;                // mm_interconnect_0:uart_so2_s1_begintransfer -> uart_so2:begintransfer
	wire  [15:0] mm_interconnect_0_uart_hmi_s1_writedata;                    // mm_interconnect_0:uart_hmi_s1_writedata -> uart_hmi:writedata
	wire   [2:0] mm_interconnect_0_uart_hmi_s1_address;                      // mm_interconnect_0:uart_hmi_s1_address -> uart_hmi:address
	wire         mm_interconnect_0_uart_hmi_s1_chipselect;                   // mm_interconnect_0:uart_hmi_s1_chipselect -> uart_hmi:chipselect
	wire         mm_interconnect_0_uart_hmi_s1_write;                        // mm_interconnect_0:uart_hmi_s1_write -> uart_hmi:write_n
	wire         mm_interconnect_0_uart_hmi_s1_read;                         // mm_interconnect_0:uart_hmi_s1_read -> uart_hmi:read_n
	wire  [15:0] mm_interconnect_0_uart_hmi_s1_readdata;                     // uart_hmi:readdata -> mm_interconnect_0:uart_hmi_s1_readdata
	wire         mm_interconnect_0_uart_hmi_s1_begintransfer;                // mm_interconnect_0:uart_hmi_s1_begintransfer -> uart_hmi:begintransfer
	wire  [15:0] mm_interconnect_0_uart_o3_s1_writedata;                     // mm_interconnect_0:uart_o3_s1_writedata -> uart_o3:writedata
	wire   [2:0] mm_interconnect_0_uart_o3_s1_address;                       // mm_interconnect_0:uart_o3_s1_address -> uart_o3:address
	wire         mm_interconnect_0_uart_o3_s1_chipselect;                    // mm_interconnect_0:uart_o3_s1_chipselect -> uart_o3:chipselect
	wire         mm_interconnect_0_uart_o3_s1_write;                         // mm_interconnect_0:uart_o3_s1_write -> uart_o3:write_n
	wire         mm_interconnect_0_uart_o3_s1_read;                          // mm_interconnect_0:uart_o3_s1_read -> uart_o3:read_n
	wire  [15:0] mm_interconnect_0_uart_o3_s1_readdata;                      // uart_o3:readdata -> mm_interconnect_0:uart_o3_s1_readdata
	wire         mm_interconnect_0_uart_o3_s1_begintransfer;                 // mm_interconnect_0:uart_o3_s1_begintransfer -> uart_o3:begintransfer
	wire   [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;         // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire  [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;        // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire         irq_mapper_receiver0_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver2_irq;                                   // key:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys:d_irq
	wire         irq_mapper_receiver1_irq;                                   // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                              // uart_no2:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver3_irq;                                   // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                          // uart_co:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver4_irq;                                   // irq_synchronizer_002:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                          // uart_sds011:irq -> irq_synchronizer_002:receiver_irq
	wire         irq_mapper_receiver5_irq;                                   // irq_synchronizer_003:sender_irq -> irq_mapper:receiver5_irq
	wire   [0:0] irq_synchronizer_003_receiver_irq;                          // uart_so2:irq -> irq_synchronizer_003:receiver_irq
	wire         irq_mapper_receiver6_irq;                                   // irq_synchronizer_004:sender_irq -> irq_mapper:receiver6_irq
	wire   [0:0] irq_synchronizer_004_receiver_irq;                          // uart_o3:irq -> irq_synchronizer_004:receiver_irq
	wire         irq_mapper_receiver7_irq;                                   // irq_synchronizer_005:sender_irq -> irq_mapper:receiver7_irq
	wire   [0:0] irq_synchronizer_005_receiver_irq;                          // uart_hmi:irq -> irq_synchronizer_005:receiver_irq
	wire         irq_mapper_receiver8_irq;                                   // irq_synchronizer_006:sender_irq -> irq_mapper:receiver8_irq
	wire   [0:0] irq_synchronizer_006_receiver_irq;                          // epcs_flash:irq -> irq_synchronizer_006:receiver_irq
	wire         rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, irq_synchronizer_005:sender_reset, irq_synchronizer_006:sender_reset, jtag_uart:rst_n, key:reset_n, mm_interconnect_0:nios2_qsys_reset_n_reset_bridge_in_reset_reset, nios2_qsys:reset_n, rst_translator:in_reset, sdram:reset_n, sysid_qsys:reset_n]
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [nios2_qsys:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_jtag_debug_module_reset_reset;                   // nios2_qsys:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [altpll:reset, epcs_flash:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, irq_synchronizer_004:receiver_reset, irq_synchronizer_005:receiver_reset, irq_synchronizer_006:receiver_reset, mm_interconnect_0:altpll_inclk_interface_reset_reset_bridge_in_reset_reset, rst_translator_001:in_reset, scl:reset_n, sda:reset_n, uart_co:reset_n, uart_hmi:reset_n, uart_no2:reset_n, uart_o3:reset_n, uart_sds011:reset_n, uart_so2:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [epcs_flash:reset_req, rst_translator_001:reset_req_in]

	DE0_NANO_QSYS_nios2_qsys nios2_qsys (
		.clk                                   (altpll_c0_clk),                                              //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                            //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                             (nios2_qsys_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                            // custom_instruction_master.readra
	);

	DE0_NANO_QSYS_sysid_qsys sysid_qsys (
		.clock    (altpll_c0_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	DE0_NANO_QSYS_jtag_uart jtag_uart (
		.clk            (altpll_c0_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	DE0_NANO_QSYS_key key (
		.clk        (altpll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver2_irq)             //                 irq.irq
	);

	DE0_NANO_QSYS_sdram sdram (
		.clk            (altpll_c0_clk),                            //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	DE0_NANO_QSYS_altpll altpll (
		.clk       (clk_clk),                                      //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),           // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_pll_slave_writedata), //                      .writedata
		.c0        (altpll_c0_clk),                                //                    c0.clk
		.c1        (altpll_sdram_clk),                             //                    c1.clk
		.areset    (altpll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (altpll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (altpll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	DE0_NANO_QSYS_scl scl (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_scl_s1_readdata),   //                    .readdata
		.out_port   (scl_export)                           // external_connection.export
	);

	DE0_NANO_QSYS_sda sda (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sda_s1_readdata),   //                    .readdata
		.bidir_port (sda_export)                           // external_connection.export
	);

	DE0_NANO_QSYS_uart_no2 uart_no2 (
		.clk           (clk_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_no2_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_no2_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_no2_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_no2_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_no2_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_no2_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_no2_s1_readdata),      //                    .readdata
		.dataavailable (),                                            //                    .dataavailable
		.readyfordata  (),                                            //                    .readyfordata
		.rxd           (uart_test_external_connection_rxd),           // external_connection.export
		.txd           (uart_test_external_connection_txd),           //                    .export
		.irq           (irq_synchronizer_receiver_irq)                //                 irq.irq
	);

	DE0_NANO_QSYS_uart_no2 uart_co (
		.clk           (clk_clk),                                    //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address       (mm_interconnect_0_uart_co_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_co_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_co_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_co_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_co_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_co_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_co_s1_readdata),      //                    .readdata
		.dataavailable (),                                           //                    .dataavailable
		.readyfordata  (),                                           //                    .readyfordata
		.rxd           (uart_co_external_connection_rxd),            // external_connection.export
		.txd           (uart_co_external_connection_txd),            //                    .export
		.irq           (irq_synchronizer_001_receiver_irq)           //                 irq.irq
	);

	DE0_NANO_QSYS_uart_no2 uart_sds011 (
		.clk           (clk_clk),                                        //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),            //               reset.reset_n
		.address       (mm_interconnect_0_uart_sds011_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_sds011_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_sds011_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_sds011_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_sds011_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_sds011_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_sds011_s1_readdata),      //                    .readdata
		.dataavailable (),                                               //                    .dataavailable
		.readyfordata  (),                                               //                    .readyfordata
		.rxd           (uart_sds011_external_connection_rxd),            // external_connection.export
		.txd           (uart_sds011_external_connection_txd),            //                    .export
		.irq           (irq_synchronizer_002_receiver_irq)               //                 irq.irq
	);

	DE0_NANO_QSYS_uart_no2 uart_so2 (
		.clk           (clk_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_so2_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_so2_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_so2_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_so2_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_so2_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_so2_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_so2_s1_readdata),      //                    .readdata
		.dataavailable (),                                            //                    .dataavailable
		.readyfordata  (),                                            //                    .readyfordata
		.rxd           (uart_so2_external_connection_rxd),            // external_connection.export
		.txd           (uart_so2_external_connection_txd),            //                    .export
		.irq           (irq_synchronizer_003_receiver_irq)            //                 irq.irq
	);

	DE0_NANO_QSYS_uart_no2 uart_o3 (
		.clk           (clk_clk),                                    //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address       (mm_interconnect_0_uart_o3_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_o3_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_o3_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_o3_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_o3_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_o3_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_o3_s1_readdata),      //                    .readdata
		.dataavailable (),                                           //                    .dataavailable
		.readyfordata  (),                                           //                    .readyfordata
		.rxd           (uart_o3_external_connection_rxd),            // external_connection.export
		.txd           (uart_o3_external_connection_txd),            //                    .export
		.irq           (irq_synchronizer_004_receiver_irq)           //                 irq.irq
	);

	DE0_NANO_QSYS_uart_hmi uart_hmi (
		.clk           (clk_clk),                                     //                 clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_hmi_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_hmi_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_hmi_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_hmi_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_hmi_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_hmi_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_hmi_s1_readdata),      //                    .readdata
		.dataavailable (),                                            //                    .dataavailable
		.readyfordata  (),                                            //                    .readyfordata
		.rxd           (uart_hmi_external_connection_rxd),            // external_connection.export
		.txd           (uart_hmi_external_connection_txd),            //                    .export
		.irq           (irq_synchronizer_005_receiver_irq)            //                 irq.irq
	);

	DE0_NANO_QSYS_epcs_flash epcs_flash (
		.clk           (clk_clk),                                                   //               clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.reset_req     (rst_controller_001_reset_out_reset_req),                    //                  .reset_req
		.address       (mm_interconnect_0_epcs_flash_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                          //                  .dataavailable
		.endofpacket   (),                                                          //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_flash_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                          //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_flash_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_synchronizer_006_receiver_irq),                         //               irq.irq
		.dclk          (epcs_flash_external_dclk),                                  //          external.export
		.sce           (epcs_flash_external_sce),                                   //                  .export
		.sdo           (epcs_flash_external_sdo),                                   //                  .export
		.data0         (epcs_flash_external_data0)                                  //                  .export
	);

	DE0_NANO_QSYS_mm_interconnect_0 mm_interconnect_0 (
		.altpll_c0_clk                                            (altpll_c0_clk),                                              //                                          altpll_c0.clk
		.clk_50_clk_clk                                           (clk_clk),                                                    //                                         clk_50_clk.clk
		.altpll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                         // altpll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_qsys_reset_n_reset_bridge_in_reset_reset           (rst_controller_reset_out_reset),                             //           nios2_qsys_reset_n_reset_bridge_in_reset.reset
		.nios2_qsys_data_master_address                           (nios2_qsys_data_master_address),                             //                             nios2_qsys_data_master.address
		.nios2_qsys_data_master_waitrequest                       (nios2_qsys_data_master_waitrequest),                         //                                                   .waitrequest
		.nios2_qsys_data_master_byteenable                        (nios2_qsys_data_master_byteenable),                          //                                                   .byteenable
		.nios2_qsys_data_master_read                              (nios2_qsys_data_master_read),                                //                                                   .read
		.nios2_qsys_data_master_readdata                          (nios2_qsys_data_master_readdata),                            //                                                   .readdata
		.nios2_qsys_data_master_readdatavalid                     (nios2_qsys_data_master_readdatavalid),                       //                                                   .readdatavalid
		.nios2_qsys_data_master_write                             (nios2_qsys_data_master_write),                               //                                                   .write
		.nios2_qsys_data_master_writedata                         (nios2_qsys_data_master_writedata),                           //                                                   .writedata
		.nios2_qsys_data_master_debugaccess                       (nios2_qsys_data_master_debugaccess),                         //                                                   .debugaccess
		.nios2_qsys_instruction_master_address                    (nios2_qsys_instruction_master_address),                      //                      nios2_qsys_instruction_master.address
		.nios2_qsys_instruction_master_waitrequest                (nios2_qsys_instruction_master_waitrequest),                  //                                                   .waitrequest
		.nios2_qsys_instruction_master_read                       (nios2_qsys_instruction_master_read),                         //                                                   .read
		.nios2_qsys_instruction_master_readdata                   (nios2_qsys_instruction_master_readdata),                     //                                                   .readdata
		.nios2_qsys_instruction_master_readdatavalid              (nios2_qsys_instruction_master_readdatavalid),                //                                                   .readdatavalid
		.altpll_pll_slave_address                                 (mm_interconnect_0_altpll_pll_slave_address),                 //                                   altpll_pll_slave.address
		.altpll_pll_slave_write                                   (mm_interconnect_0_altpll_pll_slave_write),                   //                                                   .write
		.altpll_pll_slave_read                                    (mm_interconnect_0_altpll_pll_slave_read),                    //                                                   .read
		.altpll_pll_slave_readdata                                (mm_interconnect_0_altpll_pll_slave_readdata),                //                                                   .readdata
		.altpll_pll_slave_writedata                               (mm_interconnect_0_altpll_pll_slave_writedata),               //                                                   .writedata
		.epcs_flash_epcs_control_port_address                     (mm_interconnect_0_epcs_flash_epcs_control_port_address),     //                       epcs_flash_epcs_control_port.address
		.epcs_flash_epcs_control_port_write                       (mm_interconnect_0_epcs_flash_epcs_control_port_write),       //                                                   .write
		.epcs_flash_epcs_control_port_read                        (mm_interconnect_0_epcs_flash_epcs_control_port_read),        //                                                   .read
		.epcs_flash_epcs_control_port_readdata                    (mm_interconnect_0_epcs_flash_epcs_control_port_readdata),    //                                                   .readdata
		.epcs_flash_epcs_control_port_writedata                   (mm_interconnect_0_epcs_flash_epcs_control_port_writedata),   //                                                   .writedata
		.epcs_flash_epcs_control_port_chipselect                  (mm_interconnect_0_epcs_flash_epcs_control_port_chipselect),  //                                                   .chipselect
		.jtag_uart_avalon_jtag_slave_address                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),      //                        jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),        //                                                   .write
		.jtag_uart_avalon_jtag_slave_read                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),         //                                                   .read
		.jtag_uart_avalon_jtag_slave_readdata                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),     //                                                   .readdata
		.jtag_uart_avalon_jtag_slave_writedata                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),    //                                                   .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),  //                                                   .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),   //                                                   .chipselect
		.key_s1_address                                           (mm_interconnect_0_key_s1_address),                           //                                             key_s1.address
		.key_s1_write                                             (mm_interconnect_0_key_s1_write),                             //                                                   .write
		.key_s1_readdata                                          (mm_interconnect_0_key_s1_readdata),                          //                                                   .readdata
		.key_s1_writedata                                         (mm_interconnect_0_key_s1_writedata),                         //                                                   .writedata
		.key_s1_chipselect                                        (mm_interconnect_0_key_s1_chipselect),                        //                                                   .chipselect
		.nios2_qsys_jtag_debug_module_address                     (mm_interconnect_0_nios2_qsys_jtag_debug_module_address),     //                       nios2_qsys_jtag_debug_module.address
		.nios2_qsys_jtag_debug_module_write                       (mm_interconnect_0_nios2_qsys_jtag_debug_module_write),       //                                                   .write
		.nios2_qsys_jtag_debug_module_read                        (mm_interconnect_0_nios2_qsys_jtag_debug_module_read),        //                                                   .read
		.nios2_qsys_jtag_debug_module_readdata                    (mm_interconnect_0_nios2_qsys_jtag_debug_module_readdata),    //                                                   .readdata
		.nios2_qsys_jtag_debug_module_writedata                   (mm_interconnect_0_nios2_qsys_jtag_debug_module_writedata),   //                                                   .writedata
		.nios2_qsys_jtag_debug_module_byteenable                  (mm_interconnect_0_nios2_qsys_jtag_debug_module_byteenable),  //                                                   .byteenable
		.nios2_qsys_jtag_debug_module_waitrequest                 (mm_interconnect_0_nios2_qsys_jtag_debug_module_waitrequest), //                                                   .waitrequest
		.nios2_qsys_jtag_debug_module_debugaccess                 (mm_interconnect_0_nios2_qsys_jtag_debug_module_debugaccess), //                                                   .debugaccess
		.scl_s1_address                                           (mm_interconnect_0_scl_s1_address),                           //                                             scl_s1.address
		.scl_s1_write                                             (mm_interconnect_0_scl_s1_write),                             //                                                   .write
		.scl_s1_readdata                                          (mm_interconnect_0_scl_s1_readdata),                          //                                                   .readdata
		.scl_s1_writedata                                         (mm_interconnect_0_scl_s1_writedata),                         //                                                   .writedata
		.scl_s1_chipselect                                        (mm_interconnect_0_scl_s1_chipselect),                        //                                                   .chipselect
		.sda_s1_address                                           (mm_interconnect_0_sda_s1_address),                           //                                             sda_s1.address
		.sda_s1_write                                             (mm_interconnect_0_sda_s1_write),                             //                                                   .write
		.sda_s1_readdata                                          (mm_interconnect_0_sda_s1_readdata),                          //                                                   .readdata
		.sda_s1_writedata                                         (mm_interconnect_0_sda_s1_writedata),                         //                                                   .writedata
		.sda_s1_chipselect                                        (mm_interconnect_0_sda_s1_chipselect),                        //                                                   .chipselect
		.sdram_s1_address                                         (mm_interconnect_0_sdram_s1_address),                         //                                           sdram_s1.address
		.sdram_s1_write                                           (mm_interconnect_0_sdram_s1_write),                           //                                                   .write
		.sdram_s1_read                                            (mm_interconnect_0_sdram_s1_read),                            //                                                   .read
		.sdram_s1_readdata                                        (mm_interconnect_0_sdram_s1_readdata),                        //                                                   .readdata
		.sdram_s1_writedata                                       (mm_interconnect_0_sdram_s1_writedata),                       //                                                   .writedata
		.sdram_s1_byteenable                                      (mm_interconnect_0_sdram_s1_byteenable),                      //                                                   .byteenable
		.sdram_s1_readdatavalid                                   (mm_interconnect_0_sdram_s1_readdatavalid),                   //                                                   .readdatavalid
		.sdram_s1_waitrequest                                     (mm_interconnect_0_sdram_s1_waitrequest),                     //                                                   .waitrequest
		.sdram_s1_chipselect                                      (mm_interconnect_0_sdram_s1_chipselect),                      //                                                   .chipselect
		.sysid_qsys_control_slave_address                         (mm_interconnect_0_sysid_qsys_control_slave_address),         //                           sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                        (mm_interconnect_0_sysid_qsys_control_slave_readdata),        //                                                   .readdata
		.uart_co_s1_address                                       (mm_interconnect_0_uart_co_s1_address),                       //                                         uart_co_s1.address
		.uart_co_s1_write                                         (mm_interconnect_0_uart_co_s1_write),                         //                                                   .write
		.uart_co_s1_read                                          (mm_interconnect_0_uart_co_s1_read),                          //                                                   .read
		.uart_co_s1_readdata                                      (mm_interconnect_0_uart_co_s1_readdata),                      //                                                   .readdata
		.uart_co_s1_writedata                                     (mm_interconnect_0_uart_co_s1_writedata),                     //                                                   .writedata
		.uart_co_s1_begintransfer                                 (mm_interconnect_0_uart_co_s1_begintransfer),                 //                                                   .begintransfer
		.uart_co_s1_chipselect                                    (mm_interconnect_0_uart_co_s1_chipselect),                    //                                                   .chipselect
		.uart_hmi_s1_address                                      (mm_interconnect_0_uart_hmi_s1_address),                      //                                        uart_hmi_s1.address
		.uart_hmi_s1_write                                        (mm_interconnect_0_uart_hmi_s1_write),                        //                                                   .write
		.uart_hmi_s1_read                                         (mm_interconnect_0_uart_hmi_s1_read),                         //                                                   .read
		.uart_hmi_s1_readdata                                     (mm_interconnect_0_uart_hmi_s1_readdata),                     //                                                   .readdata
		.uart_hmi_s1_writedata                                    (mm_interconnect_0_uart_hmi_s1_writedata),                    //                                                   .writedata
		.uart_hmi_s1_begintransfer                                (mm_interconnect_0_uart_hmi_s1_begintransfer),                //                                                   .begintransfer
		.uart_hmi_s1_chipselect                                   (mm_interconnect_0_uart_hmi_s1_chipselect),                   //                                                   .chipselect
		.uart_no2_s1_address                                      (mm_interconnect_0_uart_no2_s1_address),                      //                                        uart_no2_s1.address
		.uart_no2_s1_write                                        (mm_interconnect_0_uart_no2_s1_write),                        //                                                   .write
		.uart_no2_s1_read                                         (mm_interconnect_0_uart_no2_s1_read),                         //                                                   .read
		.uart_no2_s1_readdata                                     (mm_interconnect_0_uart_no2_s1_readdata),                     //                                                   .readdata
		.uart_no2_s1_writedata                                    (mm_interconnect_0_uart_no2_s1_writedata),                    //                                                   .writedata
		.uart_no2_s1_begintransfer                                (mm_interconnect_0_uart_no2_s1_begintransfer),                //                                                   .begintransfer
		.uart_no2_s1_chipselect                                   (mm_interconnect_0_uart_no2_s1_chipselect),                   //                                                   .chipselect
		.uart_o3_s1_address                                       (mm_interconnect_0_uart_o3_s1_address),                       //                                         uart_o3_s1.address
		.uart_o3_s1_write                                         (mm_interconnect_0_uart_o3_s1_write),                         //                                                   .write
		.uart_o3_s1_read                                          (mm_interconnect_0_uart_o3_s1_read),                          //                                                   .read
		.uart_o3_s1_readdata                                      (mm_interconnect_0_uart_o3_s1_readdata),                      //                                                   .readdata
		.uart_o3_s1_writedata                                     (mm_interconnect_0_uart_o3_s1_writedata),                     //                                                   .writedata
		.uart_o3_s1_begintransfer                                 (mm_interconnect_0_uart_o3_s1_begintransfer),                 //                                                   .begintransfer
		.uart_o3_s1_chipselect                                    (mm_interconnect_0_uart_o3_s1_chipselect),                    //                                                   .chipselect
		.uart_sds011_s1_address                                   (mm_interconnect_0_uart_sds011_s1_address),                   //                                     uart_sds011_s1.address
		.uart_sds011_s1_write                                     (mm_interconnect_0_uart_sds011_s1_write),                     //                                                   .write
		.uart_sds011_s1_read                                      (mm_interconnect_0_uart_sds011_s1_read),                      //                                                   .read
		.uart_sds011_s1_readdata                                  (mm_interconnect_0_uart_sds011_s1_readdata),                  //                                                   .readdata
		.uart_sds011_s1_writedata                                 (mm_interconnect_0_uart_sds011_s1_writedata),                 //                                                   .writedata
		.uart_sds011_s1_begintransfer                             (mm_interconnect_0_uart_sds011_s1_begintransfer),             //                                                   .begintransfer
		.uart_sds011_s1_chipselect                                (mm_interconnect_0_uart_sds011_s1_chipselect),                //                                                   .chipselect
		.uart_so2_s1_address                                      (mm_interconnect_0_uart_so2_s1_address),                      //                                        uart_so2_s1.address
		.uart_so2_s1_write                                        (mm_interconnect_0_uart_so2_s1_write),                        //                                                   .write
		.uart_so2_s1_read                                         (mm_interconnect_0_uart_so2_s1_read),                         //                                                   .read
		.uart_so2_s1_readdata                                     (mm_interconnect_0_uart_so2_s1_readdata),                     //                                                   .readdata
		.uart_so2_s1_writedata                                    (mm_interconnect_0_uart_so2_s1_writedata),                    //                                                   .writedata
		.uart_so2_s1_begintransfer                                (mm_interconnect_0_uart_so2_s1_begintransfer),                //                                                   .begintransfer
		.uart_so2_s1_chipselect                                   (mm_interconnect_0_uart_so2_s1_chipselect)                    //                                                   .chipselect
	);

	DE0_NANO_QSYS_irq_mapper irq_mapper (
		.clk           (altpll_c0_clk),                  //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),       // receiver8.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver5_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver6_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_005 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_005_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver7_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_006 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (altpll_c0_clk),                      //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_006_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver8_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (altpll_c0_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),           // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),       //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                           // reset_in0.reset
		.reset_in1      (nios2_qsys_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),       // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req),   //          .reset_req
		.reset_req_in0  (1'b0),                                     // (terminated)
		.reset_req_in1  (1'b0),                                     // (terminated)
		.reset_in2      (1'b0),                                     // (terminated)
		.reset_req_in2  (1'b0),                                     // (terminated)
		.reset_in3      (1'b0),                                     // (terminated)
		.reset_req_in3  (1'b0),                                     // (terminated)
		.reset_in4      (1'b0),                                     // (terminated)
		.reset_req_in4  (1'b0),                                     // (terminated)
		.reset_in5      (1'b0),                                     // (terminated)
		.reset_req_in5  (1'b0),                                     // (terminated)
		.reset_in6      (1'b0),                                     // (terminated)
		.reset_req_in6  (1'b0),                                     // (terminated)
		.reset_in7      (1'b0),                                     // (terminated)
		.reset_req_in7  (1'b0),                                     // (terminated)
		.reset_in8      (1'b0),                                     // (terminated)
		.reset_req_in8  (1'b0),                                     // (terminated)
		.reset_in9      (1'b0),                                     // (terminated)
		.reset_req_in9  (1'b0),                                     // (terminated)
		.reset_in10     (1'b0),                                     // (terminated)
		.reset_req_in10 (1'b0),                                     // (terminated)
		.reset_in11     (1'b0),                                     // (terminated)
		.reset_req_in11 (1'b0),                                     // (terminated)
		.reset_in12     (1'b0),                                     // (terminated)
		.reset_req_in12 (1'b0),                                     // (terminated)
		.reset_in13     (1'b0),                                     // (terminated)
		.reset_req_in13 (1'b0),                                     // (terminated)
		.reset_in14     (1'b0),                                     // (terminated)
		.reset_req_in14 (1'b0),                                     // (terminated)
		.reset_in15     (1'b0),                                     // (terminated)
		.reset_req_in15 (1'b0)                                      // (terminated)
	);

endmodule
